netcdf domain {
dimensions:
	x = 8 ;
	ensemble = 100 ;
variables:
	double mask(x) ;
		mask:_FillValue = -9999999. ;
	double lon(x) ;
		lon:_FillValue = -9999999. ;
	double lat(x) ;
		lat:_FillValue = -9999999. ;
	double z(x) ;
		z:_FillValue = -9999999. ;
	double part(x) ;
		part:_FillValue = -9999999. ;
	double ens(ensemble, x) ;
		ens:_FillValue = -9999999. ;
data:

 mask = 1, 1, 1, 1, 1, 1, 1, 1 ;

 lon = 1, 2, 3, 4, 5, 6, 7, 8 ;

 lat = 0, 0, 0, 0, 0, 0, 0, 0 ;

 z = 0, 0, 0, 0, 0, 0, 0, 0 ;

 part = 1, 2, 3, 4, 5, 6, 7, 8 ;

 ens =
  0.999047601928503, 1.99614220150828, 2.996428236942, 3.99156187019496, 
    4.99340568573154, 5.99861537762147, 7.01165283436256, 8.00879231347194,
  1.02350577627479, 2.00128524404712, 2.99777380411991, 3.99794568711331, 
    5.00008254877763, 6.00213723473289, 6.99726993654645, 8.00547521507156,
  1.001618587129, 1.98311896133707, 3.00487657179956, 4.00186072565143, 
    5.01582199523653, 6.00713210512924, 6.99356045389458, 8.01028218449801,
  0.993478261014915, 1.99751392173562, 2.9983082372262, 3.99535986373158, 
    5.00871523298224, 5.99491259078779, 7.00235825080396, 8.00414336405539,
  1.00835690232354, 2.01846026796573, 3.00768294857944, 3.98401109924176, 
    5.00903150288733, 6.00634138562197, 7.01517814513081, 7.99945297615412,
  1.01059748158465, 1.98835594582869, 2.9995857770166, 3.9842199444709, 
    4.9878681733941, 5.99559549324555, 7.00598607051757, 8.00847605710966,
  1.00408259225067, 1.99339179048388, 3.0057195194427, 3.99137968709225, 
    5.01149681949326, 5.98832313889525, 6.99616708339162, 8.0139001937879,
  0.980563002398504, 2.00776940621218, 3.00785043225563, 4.01123219029445, 
    5.00077931064283, 5.98305459947907, 7.00855829102211, 7.98609508597256,
  1.00858846120473, 2.00755021773058, 2.99309500710671, 4.00787459409974, 
    5.00449348767489, 6.00029669557188, 7.00465125996866, 7.99434204952393,
  1.01053631927605, 1.99145747463208, 2.98743590005122, 3.98940907184449, 
    5.00468258491803, 5.99201234474884, 7.00033335879696, 7.99469316633522,
  0.989955431474634, 2.0074088706874, 2.99862281892051, 3.99948536658867, 
    5.00387626964202, 5.99468440173788, 7.01121893249295, 7.99421111753198,
  1.01079185570858, 1.99042986808248, 2.98565876269822, 3.99891993012416, 
    5.00932362445575, 6.0056443985639, 7.00036006002472, 7.99137511452439,
  1.01184683935112, 1.99858263980388, 2.98178326394292, 3.9875029954515, 
    4.99109888991187, 5.99651716090605, 6.99267851656255, 8.00287887546247,
  1.00933715565649, 2.00286731057978, 3.00117096778405, 4.01283375966637, 
    4.99133034420431, 5.99795454436724, 7.02206012890168, 7.99380953421188,
  1.00060083469236, 1.98768422341535, 3.00797450816851, 3.98879951053073, 
    4.99571583206906, 5.98966720762472, 7.00549457517282, 8.00089072795223,
  1.00889032341285, 1.99357305090555, 3.00859750950395, 3.99277938542955, 
    4.99498433138672, 6.00993304585009, 6.99175197468784, 8.00281016889956,
  0.994701905879332, 2.01066789555686, 3.01235826054257, 4.00878710719559, 
    4.99784961967877, 6.01778145769783, 6.99308247675426, 8.00618953565134,
  0.997915157958571, 2.01337986029595, 2.99312597347906, 4.00330501702352, 
    5.01599747676594, 6.00386769921639, 7.00046330022393, 7.9959512155316,
  1.00631741558559, 1.99064123789199, 2.99131648286157, 3.99888762266248, 
    4.99369746852404, 6.00225034330985, 6.99741713879831, 8.00094919707424,
  0.98436564885708, 2.00704831110218, 3.01854262414531, 3.99785298081454, 
    5.0035855061735, 6.00283626806292, 6.99329745982573, 7.99159011650591,
  0.981600455884945, 2.00911989930108, 2.9910031093717, 4.00725012026457, 
    4.99498219957788, 5.99859279320123, 6.99607361900037, 8.00239357505982,
  1.00111243497746, 2.0171403915005, 2.9930193492702, 4.00091019159519, 
    4.99008952793819, 6.01895603700638, 7.00082900626228, 8.01371120471461,
  0.998071832785806, 1.99035606032583, 2.99525128521181, 4.02203173182934, 
    4.9953313321098, 5.99953993424847, 6.98856876754327, 8.00605617903838,
  1.01288567419716, 2.00200483117721, 3.01053579713386, 4.0054642649604, 
    5.00961375776425, 6.00531583024696, 6.99340956258639, 7.9881748348045,
  0.982769246623957, 1.98181928363377, 3.01737746604211, 3.99090170128585, 
    5.01477807994497, 6.01420804233871, 6.9943786917458, 7.99944556355767,
  1.01057709830109, 2.00386975162268, 3.02130784347177, 3.9924632631394, 
    4.99258851175048, 6.00559776811594, 6.99494693461309, 8.00949069405229,
  0.991365052182689, 1.99299454296208, 3.00687621785109, 3.99503753843618, 
    5.00404989456703, 5.98704968847929, 7.01219104509483, 7.99958949829951,
  1.00543184563347, 2.01239939640451, 3.00390726621327, 4.00742335088069, 
    5.00798954377034, 6.00887536936466, 6.99817699038557, 7.99909735132966,
  0.983576949026267, 1.98552870265034, 2.99654906456046, 3.98794667048006, 
    4.98829535000806, 5.98055822991748, 7.00239958007189, 7.99921646004229,
  1.00083533654945, 2.01528763277176, 2.99565151486764, 4.00509987385647, 
    4.99051149326654, 5.99181966916692, 6.98547649359312, 8.00729984894745,
  1.01766543877563, 1.98858960529654, 3.00582974902163, 3.98709426643498, 
    4.99642404518276, 5.98288090908172, 7.00794330036141, 8.01897587381155,
  0.9953097703631, 1.99188824643544, 3.01877606729158, 4.0031792917581, 
    4.99477105766375, 5.99263015363901, 6.98548493747733, 8.01444159626108,
  1.01326220376751, 1.98792368579052, 2.99823698305835, 4.00290914606682, 
    5.01814399259601, 5.9935001056332, 7.00325672950311, 8.01591334053279,
  1.00289637753057, 1.99596206891252, 3.02573119131711, 4.01640722441276, 
    4.98522645632521, 6.01013873338098, 7.00278256573561, 8.01613950886828,
  1.01327010263493, 1.99126916075061, 2.99144395412163, 3.97941752956032, 
    4.99083265000435, 5.99302943682451, 7.00992367968111, 8.00532545501859,
  1.00137349475958, 1.98534024421087, 3.0021957413361, 3.97511872721489, 
    5.00741482544477, 5.98911101589451, 6.98505732214197, 8.00384105078909,
  1.01857335220487, 2.01263270175779, 3.00923837884145, 3.99208097273321, 
    4.97922925734402, 6.0033109394333, 7.00872341618721, 8.00084289814631,
  1.00329804935814, 1.99539436990006, 3.0040514174286, 3.99277008893112, 
    4.99276943381851, 5.99965321086435, 6.98760323801862, 7.99192906924969,
  1.01710981660398, 1.99387910855076, 3.00695234206287, 3.99699373730694, 
    4.99924604454965, 5.99730260337678, 6.99494916274822, 7.99806901533761,
  1.00393433090998, 1.98393255266456, 2.99826970756564, 4.01010679258012, 
    4.98886638223957, 5.99649069019278, 6.99657503018055, 8.00536266500686,
  0.995202972624915, 1.99065623358832, 2.99596652253148, 4.01008188266557, 
    5.00939482848708, 6.01454993069963, 6.9902798201742, 8.00050376975829,
  1.00597365016861, 2.01197315833529, 3.00685473457571, 3.99375276715956, 
    5.00576611034125, 6.00184657208375, 7.00200904860027, 8.00094448263691,
  0.992829192548887, 1.98466037189926, 2.99925445086351, 3.99465981327734, 
    5.00631685849919, 5.98698066610407, 7.01580114032557, 8.01033524277315,
  0.984772063464235, 2.01274029989166, 3.00157968539697, 4.00692516967317, 
    5.00023023361364, 5.9881254736981, 7.01020784227602, 7.99940371030265,
  1.00403899581521, 1.99493075808274, 2.99471903794713, 3.99748764723826, 
    4.992029581285, 6.00258865950448, 7.00990805391147, 8.00070711806468,
  1.00661614722811, 2.00762637073762, 2.98499652394911, 3.99826979065242, 
    5.00612560199195, 6.01682058682387, 7.01140417972307, 7.99202827999428,
  0.994891768579635, 1.99043774623892, 2.98137757227319, 4.00323240132049, 
    5.00309972785786, 6.00648310969267, 7.01039830012946, 7.99076592953744,
  0.991910345475735, 1.99439494099021, 2.98848708390532, 3.99408722969834, 
    4.99967345769203, 6.00360847294775, 6.9802056175511, 7.99825343547325,
  0.999304390797978, 1.99722793561717, 2.99619104764327, 3.99316055023335, 
    4.99269438848221, 5.99577807999786, 6.98963662587983, 7.99537836917104,
  1.01779725860756, 2.01064018812579, 3.00322878604189, 3.99744849697078, 
    5.00781571885384, 5.98758892867928, 6.99016797793238, 7.99789473580354,
  0.996686162016731, 2.00536777815211, 3.00835034239773, 4.00208511562354, 
    4.98682067983078, 6.00528666869344, 7.00568073291202, 8.01410804281344,
  0.993334816147398, 2.01062174928583, 3.00312636824528, 3.99716117540522, 
    5.02025330007872, 5.99549091609286, 6.99119282460333, 7.98966785683658,
  1.01060572005477, 1.98341211796651, 2.99840681920242, 3.99227069134202, 
    5.00696471852097, 5.98797246088479, 7.0082900412188, 8.00814080330783,
  1.00909295744026, 1.98473189538115, 2.99732487728787, 3.9988335377779, 
    4.99734420907001, 6.00525451629777, 6.99693036305377, 7.99607150320662,
  1.00702652706946, 1.99678941978823, 3.00698434583352, 3.99863485636441, 
    4.99919105671875, 5.99226699265952, 6.9947023246101, 8.01183097876213,
  0.992007844084062, 1.99628459026905, 2.99309559563312, 3.99855235596067, 
    4.99864314662266, 6.00468359062012, 7.01018664146294, 8.00629496844337,
  0.9983480097921, 1.99171095395824, 2.9954035756545, 3.98785695934217, 
    5.0118799354957, 5.98798186724163, 6.99256276117349, 8.00289151150141,
  1.00408348745562, 2.00803553384781, 3.01700362205806, 4.01118640125013, 
    4.98873705680739, 6.01776272374844, 6.98541975455429, 8.01366787619622,
  0.994724667645564, 2.00268754620769, 3.01270566283219, 4.00284638921916, 
    5.00646305512089, 5.98301784178014, 7.00737430740259, 7.9972658827896,
  1.0166241736466, 1.99486846907078, 3.00160681923601, 4.00710301365618, 
    5.02783634256292, 5.98504045843177, 7.00532437890565, 8.00045337437893,
  0.990888236013769, 2.01567638826935, 3.00255137011301, 3.98298655810597, 
    4.99484751449337, 5.99065734214325, 7.00267507952566, 8.0047519079638,
  0.987622822689517, 1.98839046890915, 2.98875577877606, 4.00627114857152, 
    5.01287814927406, 5.98841992514714, 6.99432899063406, 7.99306803218696,
  0.998044355560549, 1.98654619453675, 2.99773541106683, 4.01105854521015, 
    5.0028449639268, 6.00279878170189, 6.99679014885321, 8.00674601939478,
  0.993987737475483, 2.00695642160346, 3.00154068387733, 3.99753722193884, 
    4.99479713446223, 6.00357055666425, 7.00519095736783, 8.00065187848958,
  1.00278963735206, 2.00586353050865, 3.00061957425641, 3.98309189241312, 
    5.01060400427876, 5.97683397827586, 6.97215389288725, 8.00166990830596,
  0.978840890093667, 2.00179403953286, 3.00307417901222, 4.00465841402655, 
    4.99838855872881, 6.01641452672582, 6.99859337958488, 7.996115693621,
  0.99733428633154, 2.00627095552451, 3.01282971509977, 3.98871557416831, 
    5.00561803242191, 5.994198901791, 7.00783972625654, 7.99511078837286,
  0.994770096537388, 1.99946480631258, 2.99539467899067, 4.01204227556194, 
    4.98151303213301, 5.98808233381643, 7.00345659537064, 8.01155807277076,
  0.982700439597973, 2.00978378441094, 3.00090442914847, 4.00372493426916, 
    4.98403600084752, 5.98471781239327, 6.99433619830556, 8.0103472990573,
  1.01532255334302, 1.98631155817266, 3.00679607181541, 4.00548940300344, 
    5.01749103211176, 6.01054610872166, 6.99586991640758, 8.02223366210431,
  1.00673992198105, 1.99107171695718, 2.99960327866043, 4.01071810154673, 
    5.00229508672218, 6.00164581867587, 7.00242708069247, 8.0067365202937,
  0.981739336086007, 1.99381401161084, 2.99388159418011, 4.01361408674719, 
    4.96769680368618, 6.00391332817282, 7.00506964105236, 8.00178250962746,
  0.987064623958822, 1.99833236596566, 2.99436114887681, 3.99674171485921, 
    4.99893038502252, 5.99948847248167, 6.97405579822209, 8.00102893700178,
  1.00011694162895, 1.99148857259165, 2.99487272315694, 4.00849364344302, 
    5.00388493115202, 5.99607922804422, 6.99172519433936, 8.0098224052622,
  0.979212152890817, 2.00237527638122, 3.00647988369423, 4.00534355899921, 
    4.98710753431222, 6.00716633680543, 6.99513089894843, 8.00736987157529,
  1.00847355922979, 1.9976037532813, 2.99318062754736, 3.9994791772141, 
    5.01056710907443, 6.02223521113587, 6.99758644828606, 8.00064030029102,
  0.997341521085403, 1.9962264068824, 3.00600566621916, 4.00525431913223, 
    4.99893656548898, 6.01430673824626, 6.98194757071601, 8.00212217712398,
  0.990122353567076, 2.00617169798912, 3.01091093691776, 4.00365752847468, 
    4.99442211723209, 5.99843374103011, 6.99700095855953, 8.00565422284661,
  1.00612116199976, 2.01418771818974, 3.02092050902839, 3.98750625553369, 
    4.99881964921485, 6.0055584805659, 7.00528585469583, 8.00163042507669,
  0.999535522934341, 1.99856662414307, 2.99446461810676, 3.98389262381627, 
    5.00256002766212, 6.01553534389288, 7.0027654787698, 8.00735735967634,
  1.00076578070151, 2.0057872118088, 2.99938922207466, 3.99879428958136, 
    5.01414495122283, 6.00896508802243, 6.99231784382078, 7.99624460285087,
  1.00279213674556, 2.00979362663884, 2.9929068612505, 4.00537757088875, 
    5.01442287317309, 5.9936854601175, 7.00310754159177, 7.9979215648147,
  1.01762498620777, 2.01894307588259, 3.0099413619835, 3.99414370836079, 
    5.0000036933941, 6.00259470390026, 6.99540114293156, 7.99325820844136,
  1.00301892477787, 2.01008824511497, 3.01342554586572, 3.99579264531967, 
    5.00292006105095, 5.99525760504255, 7.02061454666384, 7.98136529489716,
  0.997260359569149, 1.9975860375969, 2.98977811796586, 4.00547210521571, 
    4.99380927637513, 5.98643316446394, 6.99473114470967, 7.98786189561727,
  1.00135966893252, 2.00590831111503, 2.99571671420118, 4.00162091424674, 
    5.00329094682377, 6.01392656466554, 6.98372623007015, 8.03143195592816,
  1.00435860504089, 2.00416450919823, 3.00641675945154, 4.00362042464249, 
    5.0056214102407, 5.99721248158067, 7.00355409412018, 7.9995992158999,
  1.01878492002691, 2.01173954116418, 2.99313628458111, 3.98652129392329, 
    5.00957777741493, 6.02086490586055, 6.99965902035666, 7.99775386014547,
  1.0046670619254, 2.00741881768927, 3.00160487137936, 3.99132900167995, 
    5.00271813617232, 5.97411725388813, 6.99673083414783, 8.00869507483011,
  1.00209951459173, 1.99211243686889, 3.01678642461184, 4.00430937522918, 
    5.00432435584904, 6.00405195197215, 7.00798750407311, 8.00407988408578,
  1.01279090270302, 2.00206147826772, 3.00367526275663, 4.01627120707199, 
    4.99281699996636, 5.99947387772254, 7.00719440290838, 8.00866667000972,
  0.997102064726803, 2.01409381424176, 3.01561038019466, 3.99505619245715, 
    5.0158987296659, 5.98755229684998, 7.00343067588461, 8.00041008982578,
  1.01264040985493, 2.00550564406743, 3.01519606104799, 3.99622592421468, 
    5.00090996564749, 6.01835155888308, 6.98970524373881, 8.00076697982055,
  1.00554829380053, 2.01214015564984, 2.98685562016554, 3.98386615316902, 
    5.00360365349678, 6.00500982302935, 7.00341097972631, 7.99603368808808,
  1.00618646830434, 1.98998711970753, 3.01552359470061, 3.99772871640628, 
    4.99722275917696, 6.00569512461962, 6.99871413506687, 7.99496025314344,
  0.998141748878061, 1.98365796489434, 3.00332612681575, 4.01546442632123, 
    5.00840271662051, 6.00767948508063, 7.00191235663105, 7.99591630962704,
  0.987136732459278, 1.99675636283649, 2.99992054617079, 4.00658161824489, 
    5.00134341210614, 5.98662624211965, 6.98662163106084, 7.99486075285495,
  1.00363171928115, 1.98982910349261, 3.00658042991652, 3.99360972298259, 
    5.00572934495076, 6.01303402115868, 7.00783805641164, 7.99505288646338,
  1.00614863389683, 2.00904198316149, 3.00250095399209, 3.99299223489708, 
    4.99292641067237, 6.0022764338421, 6.98877705474282, 7.99889607664686,
  1.01250730582404, 2.012418980469, 3.00080536274528, 4.00719342236996, 
    4.99592866871937, 6.00538155815713, 6.98724909111248, 7.99247132816759 ;
}
